package shared_pkg;
parameter FIFO_DEPTH = 8;
parameter FIFO_WIDTH = 16;
endpackage